module mux_de_control(input [7:0] CONTROL,
                	input 		CLK,
                	input 		ENABLE,
                	input 		DIR,
			input [1:0] MODO,
			input 		S_IN,
			output reg 	S_OUT,
                        output reg [3:0] Q);
  

 
endmodule


	  
  

 



	
